-------------------------------------------
-- VHDL implementation of mu0 processor  --
-- Top level                             --
-- Ben Howes 2011                        --
-------------------------------------------
