-------------------------------------------
-- VHDL implementation of mu0 processor  --
-- Test Bench                            --
-- Ben Howes 2011                        --
-------------------------------------------
